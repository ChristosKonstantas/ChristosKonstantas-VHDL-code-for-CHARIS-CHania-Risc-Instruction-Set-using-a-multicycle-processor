--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   21:24:31 05/01/2020
-- Design Name:   
-- Module Name:   C:/Organwsi workspace/dikomou/SOURCES/ergasia1/Fetch_Ubit_TB.vhd
-- Project Name:  ergasia1
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Fetch_Unit
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY Fetch_Ubit_TB IS
END Fetch_Ubit_TB;
 
ARCHITECTURE behavior OF Fetch_Ubit_TB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Fetch_Unit
    PORT(
         PC_Immed : IN  std_logic_vector(31 downto 0);
         Instruction : OUT  std_logic_vector(31 downto 0);
         Reset : IN  std_logic;
         Clk : IN  std_logic;
         PC_LdEn : IN  std_logic;
         PC_sel : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal PC_Immed : std_logic_vector(31 downto 0) := (others => '0');
   signal Reset : std_logic := '0';
   signal Clk : std_logic := '0';
   signal PC_LdEn : std_logic := '0';
   signal PC_sel : std_logic := '0';

 	--Outputs
   signal Instruction : std_logic_vector(31 downto 0);

   -- Clock period definitions
   constant Clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Fetch_Unit PORT MAP (
          PC_Immed => PC_Immed,
          Instruction => Instruction,
          Reset => Reset,
          Clk => Clk,
          PC_LdEn => PC_LdEn,
          PC_sel => PC_sel
        );

   -- Clock process definitions
   Clk_process :process
   begin
		Clk <= '0';
		wait for Clk_period/2;
		Clk <= '1';
		wait for Clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      
		
		
    PC_Immed <= "00000000000000000000000000000001";
    Reset<='1';
    PC_LdEn<='0';
    PC_sel<='1';
      wait for Clk_period*10;
		
		PC_Immed <= "00000000000000000000000000000001";
    Reset<='0';
    PC_LdEn<='0';
    PC_sel<='1';
      wait for Clk_period*10;
		
		PC_Immed <= "00000000000000000000000000000011";
    Reset<='0';
    PC_LdEn<='0';
    PC_sel<='0';
      wait for Clk_period*10;


	PC_Immed <= "00000000000000000000000000000011";
    Reset<='0';
    PC_LdEn<='0';
    PC_sel<='0';
      wait for Clk_period*10;
		
		PC_Immed <= "00000000000000000000000000000111";
    Reset<='0';
    PC_LdEn<='0';
    PC_sel<='1';
      wait for Clk_period*10;
		
		
		PC_Immed <= "00000000000000000000000000001111";
    Reset<='0';
    PC_LdEn<='0';
    PC_sel<='0';
      wait for Clk_period*10;
      -- insert stimulus here 

      wait;
   end process;

END;
