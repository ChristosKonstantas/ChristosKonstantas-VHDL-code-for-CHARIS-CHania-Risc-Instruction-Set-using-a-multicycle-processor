
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity MEM is
end MEM;

architecture Behavioral of MEM is

begin


end Behavioral;

